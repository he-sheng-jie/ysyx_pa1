module IDU(
    input [31:0] inst,
    output [4:0] rd,
    output [4:0] rs1,
    output [4:0] rs2,
    output [31:0] imm_i,
    output [31:0] imm_u,
    output [31:0] imm_s,
    output [31:0] imm_b,
    output [31:0] imm_j,
    output [6:0] opcode,
    output [2:0] funct3,
    output [6:0] funct7
);
    assign opcode = inst[6:0];

    assign rd = inst[11:7];
    assign rs1 = inst[19:15];
    assign rs2 = inst[24:20];

    assign imm_i = { {20{inst[31]}}, inst[31:20]};
    assign imm_s = {{20{inst[31]}},inst[31:25],inst[11:7]};
    assign imm_u = {inst[31:12],12'b0};
    assign imm_b = {{20{inst[31]}},inst[7],inst[30:25],inst[11:8],1'b0};
    assign imm_j = {{11{inst[31]}},inst[31],inst[19:12],inst[20],inst[30:21],1'b0};

    assign funct3 = inst[14:12];
    assign funct7 = inst[31:25];
endmodule

