module RegisterFile #(ADDR_WIDTH = 5, DATA_WIDTH = 32) (
  input clk,
  input [DATA_WIDTH-1:0] wdata,
  input [ADDR_WIDTH-1:0] waddr,
  input wen,
  input [ADDR_WIDTH-1:0] raddr1,
  input [ADDR_WIDTH-1:0] raddr2,
  output [DATA_WIDTH-1:0] rdata1,
  output [DATA_WIDTH-1:0] rdata2,
  output [DATA_WIDTH-1:0] debug_rf [0 : 2**ADDR_WIDTH-1] 
);

  reg [DATA_WIDTH-1:0] rf [0:2**ADDR_WIDTH-1];

  initial rf[0] = 0;

  always @(posedge clk) begin
    if (wen) rf[waddr] <= wdata;  
  end

  assign rdata1 = raddr1 == 0 ? 0 : rf[raddr1];
  assign rdata2 = raddr2 == 0 ? 0 : rf[raddr2];
  assign debug_rf = rf;  

endmodule